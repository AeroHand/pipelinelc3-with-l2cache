library verilog;
use verilog.vl_types.all;
entity comp_sv_unit is
end comp_sv_unit;
